`define WidthAddr 32
