module pc_reg(
	input clk,
	input rst,
	output reg[`WidthAddr-1:0] pc,
	output reg ce
);
	


